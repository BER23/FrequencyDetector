library IEEE;
use IEEE.STD_LOGIC_1164.all;

package sdft_constant_lut is

subtype lutout is std_logic_vector (31 downto 0);
type lut is array (natural range 0 to 511) of lutout;



constant re_lut : lut :=(
	"00000000000000001111111111111010",
	"00000000000000001111111111101100",
	"00000000000000001111111111010011",
	"00000000000000001111111110110000",
	"00000000000000001111111110000100",
	"00000000000000001111111101001110",
	"00000000000000001111111100001110",
	"00000000000000001111111011000100",
	"00000000000000001111111001110000",
	"00000000000000001111111000010010",
	"00000000000000001111110110101011",
	"00000000000000001111110100111010",
	"00000000000000001111110010111111",
	"00000000000000001111110000111011",
	"00000000000000001111101110101100",
	"00000000000000001111101100010100",
	"00000000000000001111101001110010",
	"00000000000000001111100111000111",
	"00000000000000001111100100010010",
	"00000000000000001111100001010011",
	"00000000000000001111011110001011",
	"00000000000000001111011010111001",
	"00000000000000001111010111011110",
	"00000000000000001111010011111001",
	"00000000000000001111010000001011",
	"00000000000000001111001100010100",
	"00000000000000001111001000010011",
	"00000000000000001111000100001000",
	"00000000000000001110111111110101",
	"00000000000000001110111011011000",
	"00000000000000001110110110110010",
	"00000000000000001110110010000011",
	"00000000000000001110101101001010",
	"00000000000000001110101000001001",
	"00000000000000001110100010111111",
	"00000000000000001110011101101011",
	"00000000000000001110011000001111",
	"00000000000000001110010010101010",
	"00000000000000001110001100111100",
	"00000000000000001110000111000101",
	"00000000000000001110000001000110",
	"00000000000000001101111010111101",
	"00000000000000001101110100101101",
	"00000000000000001101101110010100",
	"00000000000000001101100111110010",
	"00000000000000001101100001001000",
	"00000000000000001101011010010101",
	"00000000000000001101010011011011",
	"00000000000000001101001100011000",
	"00000000000000001101000101001101",
	"00000000000000001100111101111010",
	"00000000000000001100110110011110",
	"00000000000000001100101110111011",
	"00000000000000001100100111010001",
	"00000000000000001100011111011110",
	"00000000000000001100010111100100",
	"00000000000000001100001111100010",
	"00000000000000001100000111011000",
	"00000000000000001011111111000111",
	"00000000000000001011110110101110",
	"00000000000000001011101110001111",
	"00000000000000001011100101101000",
	"00000000000000001011011100111010",
	"00000000000000001011010100000100",
	"00000000000000001011001011001000",
	"00000000000000001011000010000101",
	"00000000000000001010111000111011",
	"00000000000000001010101111101011",
	"00000000000000001010100110010100",
	"00000000000000001010011100110110",
	"00000000000000001010010011010010",
	"00000000000000001010001001100111",
	"00000000000000001001111111110110",
	"00000000000000001001110101111111",
	"00000000000000001001101100000010",
	"00000000000000001001100001111111",
	"00000000000000001001010111110110",
	"00000000000000001001001101101000",
	"00000000000000001001000011010011",
	"00000000000000001000111000111001",
	"00000000000000001000101110011010",
	"00000000000000001000100011110101",
	"00000000000000001000011001001011",
	"00000000000000001000001110011100",
	"00000000000000001000000011101000",
	"00000000000000000111111000101110",
	"00000000000000000111101101110000",
	"00000000000000000111100010101101",
	"00000000000000000111010111100110",
	"00000000000000000111001100011001",
	"00000000000000000111000001001001",
	"00000000000000000110110101110100",
	"00000000000000000110101010011011",
	"00000000000000000110011110111110",
	"00000000000000000110010011011100",
	"00000000000000000110000111110111",
	"00000000000000000101111100001110",
	"00000000000000000101110000100010",
	"00000000000000000101100100110010",
	"00000000000000000101011000111110",
	"00000000000000000101001101000111",
	"00000000000000000101000001001101",
	"00000000000000000100110101010000",
	"00000000000000000100101001010000",
	"00000000000000000100011101001101",
	"00000000000000000100010001000111",
	"00000000000000000100000100111111",
	"00000000000000000011111000110100",
	"00000000000000000011101100100110",
	"00000000000000000011100000010111",
	"00000000000000000011010100000101",
	"00000000000000000011000111110001",
	"00000000000000000010111011011100",
	"00000000000000000010101111000100",
	"00000000000000000010100010101011",
	"00000000000000000010010110010000",
	"00000000000000000010001001110100",
	"00000000000000000001111101010110",
	"00000000000000000001110000110111",
	"00000000000000000001100100011000",
	"00000000000000000001010111110111",
	"00000000000000000001001011010101",
	"00000000000000000000111110110011",
	"00000000000000000000110010010000",
	"00000000000000000000100101101100",
	"00000000000000000000011001001000",
	"00000000000000000000001100100100",
	"00000000000000000000000000000000",
	"11111111111111111111110011011100",
	"11111111111111111111100110111000",
	"11111111111111111111011010010100",
	"11111111111111111111001101110000",
	"11111111111111111111000001001101",
	"11111111111111111110110100101011",
	"11111111111111111110101000001001",
	"11111111111111111110011011101000",
	"11111111111111111110001111001001",
	"11111111111111111110000010101010",
	"11111111111111111101110110001100",
	"11111111111111111101101001110000",
	"11111111111111111101011101010101",
	"11111111111111111101010000111100",
	"11111111111111111101000100100100",
	"11111111111111111100111000001111",
	"11111111111111111100101011111011",
	"11111111111111111100011111101001",
	"11111111111111111100010011011010",
	"11111111111111111100000111001100",
	"11111111111111111011111011000001",
	"11111111111111111011101110111001",
	"11111111111111111011100010110011",
	"11111111111111111011010110110000",
	"11111111111111111011001010110000",
	"11111111111111111010111110110011",
	"11111111111111111010110010111001",
	"11111111111111111010100111000010",
	"11111111111111111010011011001110",
	"11111111111111111010001111011110",
	"11111111111111111010000011110010",
	"11111111111111111001111000001001",
	"11111111111111111001101100100100",
	"11111111111111111001100001000010",
	"11111111111111111001010101100101",
	"11111111111111111001001010001100",
	"11111111111111111000111110110111",
	"11111111111111111000110011100111",
	"11111111111111111000101000011010",
	"11111111111111111000011101010011",
	"11111111111111111000010010010000",
	"11111111111111111000000111010010",
	"11111111111111110111111100011000",
	"11111111111111110111110001100100",
	"11111111111111110111100110110101",
	"11111111111111110111011100001011",
	"11111111111111110111010001100110",
	"11111111111111110111000111000111",
	"11111111111111110110111100101101",
	"11111111111111110110110010011000",
	"11111111111111110110101000001010",
	"11111111111111110110011110000001",
	"11111111111111110110010011111110",
	"11111111111111110110001010000001",
	"11111111111111110110000000001010",
	"11111111111111110101110110011001",
	"11111111111111110101101100101110",
	"11111111111111110101100011001010",
	"11111111111111110101011001101100",
	"11111111111111110101010000010101",
	"11111111111111110101000111000101",
	"11111111111111110100111101111011",
	"11111111111111110100110100111000",
	"11111111111111110100101011111100",
	"11111111111111110100100011000110",
	"11111111111111110100011010011000",
	"11111111111111110100010001110001",
	"11111111111111110100001001010010",
	"11111111111111110100000000111001",
	"11111111111111110011111000101000",
	"11111111111111110011110000011110",
	"11111111111111110011101000011100",
	"11111111111111110011100000100010",
	"11111111111111110011011000101111",
	"11111111111111110011010001000101",
	"11111111111111110011001001100010",
	"11111111111111110011000010000110",
	"11111111111111110010111010110011",
	"11111111111111110010110011101000",
	"11111111111111110010101100100101",
	"11111111111111110010100101101011",
	"11111111111111110010011110111000",
	"11111111111111110010011000001110",
	"11111111111111110010010001101100",
	"11111111111111110010001011010011",
	"11111111111111110010000101000011",
	"11111111111111110001111110111010",
	"11111111111111110001111000111011",
	"11111111111111110001110011000100",
	"11111111111111110001101101010110",
	"11111111111111110001100111110001",
	"11111111111111110001100010010101",
	"11111111111111110001011101000001",
	"11111111111111110001010111110111",
	"11111111111111110001010010110110",
	"11111111111111110001001101111101",
	"11111111111111110001001001001110",
	"11111111111111110001000100101000",
	"11111111111111110001000000001011",
	"11111111111111110000111011111000",
	"11111111111111110000110111101101",
	"11111111111111110000110011101100",
	"11111111111111110000101111110101",
	"11111111111111110000101100000111",
	"11111111111111110000101000100010",
	"11111111111111110000100101000111",
	"11111111111111110000100001110101",
	"11111111111111110000011110101101",
	"11111111111111110000011011101110",
	"11111111111111110000011000111001",
	"11111111111111110000010110001110",
	"11111111111111110000010011101100",
	"11111111111111110000010001010100",
	"11111111111111110000001111000101",
	"11111111111111110000001101000001",
	"11111111111111110000001011000110",
	"11111111111111110000001001010101",
	"11111111111111110000000111101110",
	"11111111111111110000000110010000",
	"11111111111111110000000100111100",
	"11111111111111110000000011110010",
	"11111111111111110000000010110010",
	"11111111111111110000000001111100",
	"11111111111111110000000001010000",
	"11111111111111110000000000101101",
	"11111111111111110000000000010100",
	"11111111111111110000000000000110",
	"11111111111111110000000000000001",
	"11111111111111110000000000000110",
	"11111111111111110000000000010100",
	"11111111111111110000000000101101",
	"11111111111111110000000001010000",
	"11111111111111110000000001111100",
	"11111111111111110000000010110010",
	"11111111111111110000000011110010",
	"11111111111111110000000100111100",
	"11111111111111110000000110010000",
	"11111111111111110000000111101110",
	"11111111111111110000001001010101",
	"11111111111111110000001011000110",
	"11111111111111110000001101000001",
	"11111111111111110000001111000101",
	"11111111111111110000010001010100",
	"11111111111111110000010011101100",
	"11111111111111110000010110001110",
	"11111111111111110000011000111001",
	"11111111111111110000011011101110",
	"11111111111111110000011110101101",
	"11111111111111110000100001110101",
	"11111111111111110000100101000111",
	"11111111111111110000101000100010",
	"11111111111111110000101100000111",
	"11111111111111110000101111110101",
	"11111111111111110000110011101100",
	"11111111111111110000110111101101",
	"11111111111111110000111011111000",
	"11111111111111110001000000001011",
	"11111111111111110001000100101000",
	"11111111111111110001001001001110",
	"11111111111111110001001101111101",
	"11111111111111110001010010110110",
	"11111111111111110001010111110111",
	"11111111111111110001011101000001",
	"11111111111111110001100010010101",
	"11111111111111110001100111110001",
	"11111111111111110001101101010110",
	"11111111111111110001110011000100",
	"11111111111111110001111000111011",
	"11111111111111110001111110111010",
	"11111111111111110010000101000011",
	"11111111111111110010001011010011",
	"11111111111111110010010001101100",
	"11111111111111110010011000001110",
	"11111111111111110010011110111000",
	"11111111111111110010100101101011",
	"11111111111111110010101100100101",
	"11111111111111110010110011101000",
	"11111111111111110010111010110011",
	"11111111111111110011000010000110",
	"11111111111111110011001001100010",
	"11111111111111110011010001000101",
	"11111111111111110011011000101111",
	"11111111111111110011100000100010",
	"11111111111111110011101000011100",
	"11111111111111110011110000011110",
	"11111111111111110011111000101000",
	"11111111111111110100000000111001",
	"11111111111111110100001001010010",
	"11111111111111110100010001110001",
	"11111111111111110100011010011000",
	"11111111111111110100100011000110",
	"11111111111111110100101011111100",
	"11111111111111110100110100111000",
	"11111111111111110100111101111011",
	"11111111111111110101000111000101",
	"11111111111111110101010000010101",
	"11111111111111110101011001101100",
	"11111111111111110101100011001010",
	"11111111111111110101101100101110",
	"11111111111111110101110110011001",
	"11111111111111110110000000001010",
	"11111111111111110110001010000001",
	"11111111111111110110010011111110",
	"11111111111111110110011110000001",
	"11111111111111110110101000001010",
	"11111111111111110110110010011000",
	"11111111111111110110111100101101",
	"11111111111111110111000111000111",
	"11111111111111110111010001100110",
	"11111111111111110111011100001011",
	"11111111111111110111100110110101",
	"11111111111111110111110001100100",
	"11111111111111110111111100011000",
	"11111111111111111000000111010010",
	"11111111111111111000010010010000",
	"11111111111111111000011101010011",
	"11111111111111111000101000011010",
	"11111111111111111000110011100111",
	"11111111111111111000111110110111",
	"11111111111111111001001010001100",
	"11111111111111111001010101100101",
	"11111111111111111001100001000010",
	"11111111111111111001101100100100",
	"11111111111111111001111000001001",
	"11111111111111111010000011110010",
	"11111111111111111010001111011110",
	"11111111111111111010011011001110",
	"11111111111111111010100111000010",
	"11111111111111111010110010111001",
	"11111111111111111010111110110011",
	"11111111111111111011001010110000",
	"11111111111111111011010110110000",
	"11111111111111111011100010110011",
	"11111111111111111011101110111001",
	"11111111111111111011111011000001",
	"11111111111111111100000111001100",
	"11111111111111111100010011011010",
	"11111111111111111100011111101001",
	"11111111111111111100101011111011",
	"11111111111111111100111000001111",
	"11111111111111111101000100100100",
	"11111111111111111101010000111100",
	"11111111111111111101011101010101",
	"11111111111111111101101001110000",
	"11111111111111111101110110001100",
	"11111111111111111110000010101010",
	"11111111111111111110001111001001",
	"11111111111111111110011011101000",
	"11111111111111111110101000001001",
	"11111111111111111110110100101011",
	"11111111111111111111000001001101",
	"11111111111111111111001101110000",
	"11111111111111111111011010010100",
	"11111111111111111111100110111000",
	"11111111111111111111110011011100",
	"00000000000000000000000000000000",
	"00000000000000000000001100100100",
	"00000000000000000000011001001000",
	"00000000000000000000100101101100",
	"00000000000000000000110010010000",
	"00000000000000000000111110110011",
	"00000000000000000001001011010101",
	"00000000000000000001010111110111",
	"00000000000000000001100100011000",
	"00000000000000000001110000110111",
	"00000000000000000001111101010110",
	"00000000000000000010001001110100",
	"00000000000000000010010110010000",
	"00000000000000000010100010101011",
	"00000000000000000010101111000100",
	"00000000000000000010111011011100",
	"00000000000000000011000111110001",
	"00000000000000000011010100000101",
	"00000000000000000011100000010111",
	"00000000000000000011101100100110",
	"00000000000000000011111000110100",
	"00000000000000000100000100111111",
	"00000000000000000100010001000111",
	"00000000000000000100011101001101",
	"00000000000000000100101001010000",
	"00000000000000000100110101010000",
	"00000000000000000101000001001101",
	"00000000000000000101001101000111",
	"00000000000000000101011000111110",
	"00000000000000000101100100110010",
	"00000000000000000101110000100010",
	"00000000000000000101111100001110",
	"00000000000000000110000111110111",
	"00000000000000000110010011011100",
	"00000000000000000110011110111110",
	"00000000000000000110101010011011",
	"00000000000000000110110101110100",
	"00000000000000000111000001001001",
	"00000000000000000111001100011001",
	"00000000000000000111010111100110",
	"00000000000000000111100010101101",
	"00000000000000000111101101110000",
	"00000000000000000111111000101110",
	"00000000000000001000000011101000",
	"00000000000000001000001110011100",
	"00000000000000001000011001001011",
	"00000000000000001000100011110101",
	"00000000000000001000101110011010",
	"00000000000000001000111000111001",
	"00000000000000001001000011010011",
	"00000000000000001001001101101000",
	"00000000000000001001010111110110",
	"00000000000000001001100001111111",
	"00000000000000001001101100000010",
	"00000000000000001001110101111111",
	"00000000000000001001111111110110",
	"00000000000000001010001001100111",
	"00000000000000001010010011010010",
	"00000000000000001010011100110110",
	"00000000000000001010100110010100",
	"00000000000000001010101111101011",
	"00000000000000001010111000111011",
	"00000000000000001011000010000101",
	"00000000000000001011001011001000",
	"00000000000000001011010100000100",
	"00000000000000001011011100111010",
	"00000000000000001011100101101000",
	"00000000000000001011101110001111",
	"00000000000000001011110110101110",
	"00000000000000001011111111000111",
	"00000000000000001100000111011000",
	"00000000000000001100001111100010",
	"00000000000000001100010111100100",
	"00000000000000001100011111011110",
	"00000000000000001100100111010001",
	"00000000000000001100101110111011",
	"00000000000000001100110110011110",
	"00000000000000001100111101111010",
	"00000000000000001101000101001101",
	"00000000000000001101001100011000",
	"00000000000000001101010011011011",
	"00000000000000001101011010010101",
	"00000000000000001101100001001000",
	"00000000000000001101100111110010",
	"00000000000000001101101110010100",
	"00000000000000001101110100101101",
	"00000000000000001101111010111101",
	"00000000000000001110000001000110",
	"00000000000000001110000111000101",
	"00000000000000001110001100111100",
	"00000000000000001110010010101010",
	"00000000000000001110011000001111",
	"00000000000000001110011101101011",
	"00000000000000001110100010111111",
	"00000000000000001110101000001001",
	"00000000000000001110101101001010",
	"00000000000000001110110010000011",
	"00000000000000001110110110110010",
	"00000000000000001110111011011000",
	"00000000000000001110111111110101",
	"00000000000000001111000100001000",
	"00000000000000001111001000010011",
	"00000000000000001111001100010100",
	"00000000000000001111010000001011",
	"00000000000000001111010011111001",
	"00000000000000001111010111011110",
	"00000000000000001111011010111001",
	"00000000000000001111011110001011",
	"00000000000000001111100001010011",
	"00000000000000001111100100010010",
	"00000000000000001111100111000111",
	"00000000000000001111101001110010",
	"00000000000000001111101100010100",
	"00000000000000001111101110101100",
	"00000000000000001111110000111011",
	"00000000000000001111110010111111",
	"00000000000000001111110100111010",
	"00000000000000001111110110101011",
	"00000000000000001111111000010010",
	"00000000000000001111111001110000",
	"00000000000000001111111011000100",
	"00000000000000001111111100001110",
	"00000000000000001111111101001110",
	"00000000000000001111111110000100",
	"00000000000000001111111110110000",
	"00000000000000001111111111010011",
	"00000000000000001111111111101100",
	"00000000000000001111111111111010",
	"00000000000000001111111111111111"
);
 
constant im_lut : lut :=( 
 	"00000000000000000000001100100100",
	"00000000000000000000011001001000",
	"00000000000000000000100101101100",
	"00000000000000000000110010010000",
	"00000000000000000000111110110011",
	"00000000000000000001001011010101",
	"00000000000000000001010111110111",
	"00000000000000000001100100011000",
	"00000000000000000001110000110111",
	"00000000000000000001111101010110",
	"00000000000000000010001001110100",
	"00000000000000000010010110010000",
	"00000000000000000010100010101011",
	"00000000000000000010101111000100",
	"00000000000000000010111011011100",
	"00000000000000000011000111110001",
	"00000000000000000011010100000101",
	"00000000000000000011100000010111",
	"00000000000000000011101100100110",
	"00000000000000000011111000110100",
	"00000000000000000100000100111111",
	"00000000000000000100010001000111",
	"00000000000000000100011101001101",
	"00000000000000000100101001010000",
	"00000000000000000100110101010000",
	"00000000000000000101000001001101",
	"00000000000000000101001101000111",
	"00000000000000000101011000111110",
	"00000000000000000101100100110010",
	"00000000000000000101110000100010",
	"00000000000000000101111100001110",
	"00000000000000000110000111110111",
	"00000000000000000110010011011100",
	"00000000000000000110011110111110",
	"00000000000000000110101010011011",
	"00000000000000000110110101110100",
	"00000000000000000111000001001001",
	"00000000000000000111001100011001",
	"00000000000000000111010111100110",
	"00000000000000000111100010101101",
	"00000000000000000111101101110000",
	"00000000000000000111111000101110",
	"00000000000000001000000011101000",
	"00000000000000001000001110011100",
	"00000000000000001000011001001011",
	"00000000000000001000100011110101",
	"00000000000000001000101110011010",
	"00000000000000001000111000111001",
	"00000000000000001001000011010011",
	"00000000000000001001001101101000",
	"00000000000000001001010111110110",
	"00000000000000001001100001111111",
	"00000000000000001001101100000010",
	"00000000000000001001110101111111",
	"00000000000000001001111111110110",
	"00000000000000001010001001100111",
	"00000000000000001010010011010010",
	"00000000000000001010011100110110",
	"00000000000000001010100110010100",
	"00000000000000001010101111101011",
	"00000000000000001010111000111011",
	"00000000000000001011000010000101",
	"00000000000000001011001011001000",
	"00000000000000001011010100000100",
	"00000000000000001011011100111010",
	"00000000000000001011100101101000",
	"00000000000000001011101110001111",
	"00000000000000001011110110101110",
	"00000000000000001011111111000111",
	"00000000000000001100000111011000",
	"00000000000000001100001111100010",
	"00000000000000001100010111100100",
	"00000000000000001100011111011110",
	"00000000000000001100100111010001",
	"00000000000000001100101110111011",
	"00000000000000001100110110011110",
	"00000000000000001100111101111010",
	"00000000000000001101000101001101",
	"00000000000000001101001100011000",
	"00000000000000001101010011011011",
	"00000000000000001101011010010101",
	"00000000000000001101100001001000",
	"00000000000000001101100111110010",
	"00000000000000001101101110010100",
	"00000000000000001101110100101101",
	"00000000000000001101111010111101",
	"00000000000000001110000001000110",
	"00000000000000001110000111000101",
	"00000000000000001110001100111100",
	"00000000000000001110010010101010",
	"00000000000000001110011000001111",
	"00000000000000001110011101101011",
	"00000000000000001110100010111111",
	"00000000000000001110101000001001",
	"00000000000000001110101101001010",
	"00000000000000001110110010000011",
	"00000000000000001110110110110010",
	"00000000000000001110111011011000",
	"00000000000000001110111111110101",
	"00000000000000001111000100001000",
	"00000000000000001111001000010011",
	"00000000000000001111001100010100",
	"00000000000000001111010000001011",
	"00000000000000001111010011111001",
	"00000000000000001111010111011110",
	"00000000000000001111011010111001",
	"00000000000000001111011110001011",
	"00000000000000001111100001010011",
	"00000000000000001111100100010010",
	"00000000000000001111100111000111",
	"00000000000000001111101001110010",
	"00000000000000001111101100010100",
	"00000000000000001111101110101100",
	"00000000000000001111110000111011",
	"00000000000000001111110010111111",
	"00000000000000001111110100111010",
	"00000000000000001111110110101011",
	"00000000000000001111111000010010",
	"00000000000000001111111001110000",
	"00000000000000001111111011000100",
	"00000000000000001111111100001110",
	"00000000000000001111111101001110",
	"00000000000000001111111110000100",
	"00000000000000001111111110110000",
	"00000000000000001111111111010011",
	"00000000000000001111111111101100",
	"00000000000000001111111111111010",
	"00000000000000001111111111111111",
	"00000000000000001111111111111010",
	"00000000000000001111111111101100",
	"00000000000000001111111111010011",
	"00000000000000001111111110110000",
	"00000000000000001111111110000100",
	"00000000000000001111111101001110",
	"00000000000000001111111100001110",
	"00000000000000001111111011000100",
	"00000000000000001111111001110000",
	"00000000000000001111111000010010",
	"00000000000000001111110110101011",
	"00000000000000001111110100111010",
	"00000000000000001111110010111111",
	"00000000000000001111110000111011",
	"00000000000000001111101110101100",
	"00000000000000001111101100010100",
	"00000000000000001111101001110010",
	"00000000000000001111100111000111",
	"00000000000000001111100100010010",
	"00000000000000001111100001010011",
	"00000000000000001111011110001011",
	"00000000000000001111011010111001",
	"00000000000000001111010111011110",
	"00000000000000001111010011111001",
	"00000000000000001111010000001011",
	"00000000000000001111001100010100",
	"00000000000000001111001000010011",
	"00000000000000001111000100001000",
	"00000000000000001110111111110101",
	"00000000000000001110111011011000",
	"00000000000000001110110110110010",
	"00000000000000001110110010000011",
	"00000000000000001110101101001010",
	"00000000000000001110101000001001",
	"00000000000000001110100010111111",
	"00000000000000001110011101101011",
	"00000000000000001110011000001111",
	"00000000000000001110010010101010",
	"00000000000000001110001100111100",
	"00000000000000001110000111000101",
	"00000000000000001110000001000110",
	"00000000000000001101111010111101",
	"00000000000000001101110100101101",
	"00000000000000001101101110010100",
	"00000000000000001101100111110010",
	"00000000000000001101100001001000",
	"00000000000000001101011010010101",
	"00000000000000001101010011011011",
	"00000000000000001101001100011000",
	"00000000000000001101000101001101",
	"00000000000000001100111101111010",
	"00000000000000001100110110011110",
	"00000000000000001100101110111011",
	"00000000000000001100100111010001",
	"00000000000000001100011111011110",
	"00000000000000001100010111100100",
	"00000000000000001100001111100010",
	"00000000000000001100000111011000",
	"00000000000000001011111111000111",
	"00000000000000001011110110101110",
	"00000000000000001011101110001111",
	"00000000000000001011100101101000",
	"00000000000000001011011100111010",
	"00000000000000001011010100000100",
	"00000000000000001011001011001000",
	"00000000000000001011000010000101",
	"00000000000000001010111000111011",
	"00000000000000001010101111101011",
	"00000000000000001010100110010100",
	"00000000000000001010011100110110",
	"00000000000000001010010011010010",
	"00000000000000001010001001100111",
	"00000000000000001001111111110110",
	"00000000000000001001110101111111",
	"00000000000000001001101100000010",
	"00000000000000001001100001111111",
	"00000000000000001001010111110110",
	"00000000000000001001001101101000",
	"00000000000000001001000011010011",
	"00000000000000001000111000111001",
	"00000000000000001000101110011010",
	"00000000000000001000100011110101",
	"00000000000000001000011001001011",
	"00000000000000001000001110011100",
	"00000000000000001000000011101000",
	"00000000000000000111111000101110",
	"00000000000000000111101101110000",
	"00000000000000000111100010101101",
	"00000000000000000111010111100110",
	"00000000000000000111001100011001",
	"00000000000000000111000001001001",
	"00000000000000000110110101110100",
	"00000000000000000110101010011011",
	"00000000000000000110011110111110",
	"00000000000000000110010011011100",
	"00000000000000000110000111110111",
	"00000000000000000101111100001110",
	"00000000000000000101110000100010",
	"00000000000000000101100100110010",
	"00000000000000000101011000111110",
	"00000000000000000101001101000111",
	"00000000000000000101000001001101",
	"00000000000000000100110101010000",
	"00000000000000000100101001010000",
	"00000000000000000100011101001101",
	"00000000000000000100010001000111",
	"00000000000000000100000100111111",
	"00000000000000000011111000110100",
	"00000000000000000011101100100110",
	"00000000000000000011100000010111",
	"00000000000000000011010100000101",
	"00000000000000000011000111110001",
	"00000000000000000010111011011100",
	"00000000000000000010101111000100",
	"00000000000000000010100010101011",
	"00000000000000000010010110010000",
	"00000000000000000010001001110100",
	"00000000000000000001111101010110",
	"00000000000000000001110000110111",
	"00000000000000000001100100011000",
	"00000000000000000001010111110111",
	"00000000000000000001001011010101",
	"00000000000000000000111110110011",
	"00000000000000000000110010010000",
	"00000000000000000000100101101100",
	"00000000000000000000011001001000",
	"00000000000000000000001100100100",
	"00000000000000000000000000000000",
	"11111111111111111111110011011100",
	"11111111111111111111100110111000",
	"11111111111111111111011010010100",
	"11111111111111111111001101110000",
	"11111111111111111111000001001101",
	"11111111111111111110110100101011",
	"11111111111111111110101000001001",
	"11111111111111111110011011101000",
	"11111111111111111110001111001001",
	"11111111111111111110000010101010",
	"11111111111111111101110110001100",
	"11111111111111111101101001110000",
	"11111111111111111101011101010101",
	"11111111111111111101010000111100",
	"11111111111111111101000100100100",
	"11111111111111111100111000001111",
	"11111111111111111100101011111011",
	"11111111111111111100011111101001",
	"11111111111111111100010011011010",
	"11111111111111111100000111001100",
	"11111111111111111011111011000001",
	"11111111111111111011101110111001",
	"11111111111111111011100010110011",
	"11111111111111111011010110110000",
	"11111111111111111011001010110000",
	"11111111111111111010111110110011",
	"11111111111111111010110010111001",
	"11111111111111111010100111000010",
	"11111111111111111010011011001110",
	"11111111111111111010001111011110",
	"11111111111111111010000011110010",
	"11111111111111111001111000001001",
	"11111111111111111001101100100100",
	"11111111111111111001100001000010",
	"11111111111111111001010101100101",
	"11111111111111111001001010001100",
	"11111111111111111000111110110111",
	"11111111111111111000110011100111",
	"11111111111111111000101000011010",
	"11111111111111111000011101010011",
	"11111111111111111000010010010000",
	"11111111111111111000000111010010",
	"11111111111111110111111100011000",
	"11111111111111110111110001100100",
	"11111111111111110111100110110101",
	"11111111111111110111011100001011",
	"11111111111111110111010001100110",
	"11111111111111110111000111000111",
	"11111111111111110110111100101101",
	"11111111111111110110110010011000",
	"11111111111111110110101000001010",
	"11111111111111110110011110000001",
	"11111111111111110110010011111110",
	"11111111111111110110001010000001",
	"11111111111111110110000000001010",
	"11111111111111110101110110011001",
	"11111111111111110101101100101110",
	"11111111111111110101100011001010",
	"11111111111111110101011001101100",
	"11111111111111110101010000010101",
	"11111111111111110101000111000101",
	"11111111111111110100111101111011",
	"11111111111111110100110100111000",
	"11111111111111110100101011111100",
	"11111111111111110100100011000110",
	"11111111111111110100011010011000",
	"11111111111111110100010001110001",
	"11111111111111110100001001010010",
	"11111111111111110100000000111001",
	"11111111111111110011111000101000",
	"11111111111111110011110000011110",
	"11111111111111110011101000011100",
	"11111111111111110011100000100010",
	"11111111111111110011011000101111",
	"11111111111111110011010001000101",
	"11111111111111110011001001100010",
	"11111111111111110011000010000110",
	"11111111111111110010111010110011",
	"11111111111111110010110011101000",
	"11111111111111110010101100100101",
	"11111111111111110010100101101011",
	"11111111111111110010011110111000",
	"11111111111111110010011000001110",
	"11111111111111110010010001101100",
	"11111111111111110010001011010011",
	"11111111111111110010000101000011",
	"11111111111111110001111110111010",
	"11111111111111110001111000111011",
	"11111111111111110001110011000100",
	"11111111111111110001101101010110",
	"11111111111111110001100111110001",
	"11111111111111110001100010010101",
	"11111111111111110001011101000001",
	"11111111111111110001010111110111",
	"11111111111111110001010010110110",
	"11111111111111110001001101111101",
	"11111111111111110001001001001110",
	"11111111111111110001000100101000",
	"11111111111111110001000000001011",
	"11111111111111110000111011111000",
	"11111111111111110000110111101101",
	"11111111111111110000110011101100",
	"11111111111111110000101111110101",
	"11111111111111110000101100000111",
	"11111111111111110000101000100010",
	"11111111111111110000100101000111",
	"11111111111111110000100001110101",
	"11111111111111110000011110101101",
	"11111111111111110000011011101110",
	"11111111111111110000011000111001",
	"11111111111111110000010110001110",
	"11111111111111110000010011101100",
	"11111111111111110000010001010100",
	"11111111111111110000001111000101",
	"11111111111111110000001101000001",
	"11111111111111110000001011000110",
	"11111111111111110000001001010101",
	"11111111111111110000000111101110",
	"11111111111111110000000110010000",
	"11111111111111110000000100111100",
	"11111111111111110000000011110010",
	"11111111111111110000000010110010",
	"11111111111111110000000001111100",
	"11111111111111110000000001010000",
	"11111111111111110000000000101101",
	"11111111111111110000000000010100",
	"11111111111111110000000000000110",
	"11111111111111110000000000000001",
	"11111111111111110000000000000110",
	"11111111111111110000000000010100",
	"11111111111111110000000000101101",
	"11111111111111110000000001010000",
	"11111111111111110000000001111100",
	"11111111111111110000000010110010",
	"11111111111111110000000011110010",
	"11111111111111110000000100111100",
	"11111111111111110000000110010000",
	"11111111111111110000000111101110",
	"11111111111111110000001001010101",
	"11111111111111110000001011000110",
	"11111111111111110000001101000001",
	"11111111111111110000001111000101",
	"11111111111111110000010001010100",
	"11111111111111110000010011101100",
	"11111111111111110000010110001110",
	"11111111111111110000011000111001",
	"11111111111111110000011011101110",
	"11111111111111110000011110101101",
	"11111111111111110000100001110101",
	"11111111111111110000100101000111",
	"11111111111111110000101000100010",
	"11111111111111110000101100000111",
	"11111111111111110000101111110101",
	"11111111111111110000110011101100",
	"11111111111111110000110111101101",
	"11111111111111110000111011111000",
	"11111111111111110001000000001011",
	"11111111111111110001000100101000",
	"11111111111111110001001001001110",
	"11111111111111110001001101111101",
	"11111111111111110001010010110110",
	"11111111111111110001010111110111",
	"11111111111111110001011101000001",
	"11111111111111110001100010010101",
	"11111111111111110001100111110001",
	"11111111111111110001101101010110",
	"11111111111111110001110011000100",
	"11111111111111110001111000111011",
	"11111111111111110001111110111010",
	"11111111111111110010000101000011",
	"11111111111111110010001011010011",
	"11111111111111110010010001101100",
	"11111111111111110010011000001110",
	"11111111111111110010011110111000",
	"11111111111111110010100101101011",
	"11111111111111110010101100100101",
	"11111111111111110010110011101000",
	"11111111111111110010111010110011",
	"11111111111111110011000010000110",
	"11111111111111110011001001100010",
	"11111111111111110011010001000101",
	"11111111111111110011011000101111",
	"11111111111111110011100000100010",
	"11111111111111110011101000011100",
	"11111111111111110011110000011110",
	"11111111111111110011111000101000",
	"11111111111111110100000000111001",
	"11111111111111110100001001010010",
	"11111111111111110100010001110001",
	"11111111111111110100011010011000",
	"11111111111111110100100011000110",
	"11111111111111110100101011111100",
	"11111111111111110100110100111000",
	"11111111111111110100111101111011",
	"11111111111111110101000111000101",
	"11111111111111110101010000010101",
	"11111111111111110101011001101100",
	"11111111111111110101100011001010",
	"11111111111111110101101100101110",
	"11111111111111110101110110011001",
	"11111111111111110110000000001010",
	"11111111111111110110001010000001",
	"11111111111111110110010011111110",
	"11111111111111110110011110000001",
	"11111111111111110110101000001010",
	"11111111111111110110110010011000",
	"11111111111111110110111100101101",
	"11111111111111110111000111000111",
	"11111111111111110111010001100110",
	"11111111111111110111011100001011",
	"11111111111111110111100110110101",
	"11111111111111110111110001100100",
	"11111111111111110111111100011000",
	"11111111111111111000000111010010",
	"11111111111111111000010010010000",
	"11111111111111111000011101010011",
	"11111111111111111000101000011010",
	"11111111111111111000110011100111",
	"11111111111111111000111110110111",
	"11111111111111111001001010001100",
	"11111111111111111001010101100101",
	"11111111111111111001100001000010",
	"11111111111111111001101100100100",
	"11111111111111111001111000001001",
	"11111111111111111010000011110010",
	"11111111111111111010001111011110",
	"11111111111111111010011011001110",
	"11111111111111111010100111000010",
	"11111111111111111010110010111001",
	"11111111111111111010111110110011",
	"11111111111111111011001010110000",
	"11111111111111111011010110110000",
	"11111111111111111011100010110011",
	"11111111111111111011101110111001",
	"11111111111111111011111011000001",
	"11111111111111111100000111001100",
	"11111111111111111100010011011010",
	"11111111111111111100011111101001",
	"11111111111111111100101011111011",
	"11111111111111111100111000001111",
	"11111111111111111101000100100100",
	"11111111111111111101010000111100",
	"11111111111111111101011101010101",
	"11111111111111111101101001110000",
	"11111111111111111101110110001100",
	"11111111111111111110000010101010",
	"11111111111111111110001111001001",
	"11111111111111111110011011101000",
	"11111111111111111110101000001001",
	"11111111111111111110110100101011",
	"11111111111111111111000001001101",
	"11111111111111111111001101110000",
	"11111111111111111111011010010100",
	"11111111111111111111100110111000",
	"11111111111111111111110011011100",
	"00000000000000000000000000000000"
 );
 
 end sdft_constant_lut;

package body sdft_constant_lut is
 
end sdft_constant_lut;
